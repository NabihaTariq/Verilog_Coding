`define locations 8
`define location_size 8